package defs;

typedef enum {
    ADD,
    SUB,
    DIV,
    MUL
} OP_T;

`include "checker.sv"
`include "generator.sv"

endpackage : defs
