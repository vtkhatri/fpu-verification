class common;

    static mailbox gen2drv = new();
    static mailbox mon2cov = new();
    static mailbox mon2che = new();
    static virtual bfm cbfm0;

endclass : common