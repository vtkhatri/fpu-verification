typedef enum {
    ADD,
    SUB,
    DIV,
    MUL
} OP_T;
