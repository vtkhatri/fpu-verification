class scoreboard;






endclass