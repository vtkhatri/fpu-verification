`timescale 1ns/100ps

`include "../duv/fpu.v"

`include "defs.sv"
`include "generator.sv"
`include "checker.sv"
// `include "scoreboard.sv"
