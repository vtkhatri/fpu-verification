class common;

    static mailbox gen2drv = new();
    static mailbox mon2sco = new();
    static virtual bfm sif;

endclass : common