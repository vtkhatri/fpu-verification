`timescale 1ns/100ps

`include "../duv/pre_norm_fmul.v"
`include "../duv/primitives.v"
`include "../duv/post_norm.v"
`include "../duv/pre_norm.v"
`include "../duv/except.v"
`include "../duv/fpu.v"

`include "defs.sv"
`include "generator.sv"
// `include "checker.sv"
// `include "scoreboard.sv"
