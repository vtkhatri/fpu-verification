typedef enum {
    ADD,
    SUB,
    MUL,
    DIV
} OP_T;
